module Not_gate(
	input wire a,
	output wire y
);

  assign y = ~a;

endmodule